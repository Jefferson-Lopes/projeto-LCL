module sistemaDeControle (SW, KEY);
	input [9:0] SW;
	input [3:0] KEY;


endmodule
